/****************************************************************************
 * pss_port.svh
 ****************************************************************************/

/**
 * Class: pss_port
 * 
 * TODO: Add class documentation
 */
class pss_port #(type interface_t) extends pss_port_base;
	interface_t					ifc;

	function new(string name, pss_graph parent);
		super.new(name, parent);
	endfunction

endclass

