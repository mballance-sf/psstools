/****************************************************************************
 * reg2axi_top.svh
 ****************************************************************************/

/**
 * Class: reg2axi_top
 * 
 * TODO: Add class documentation
 */
class reg2axi_top;

	function new();

	endfunction


endclass

