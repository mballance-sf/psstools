/****************************************************************************
 * pss_stdlib_pkg.sv
 ****************************************************************************/

/**
 * Package: pss_stdlib_pkg
 * 
 * TODO: Add package documentation
 */
package pss_stdlib_pkg;
	`include "pss_graph.svh"
	`include "pss_port_base.svh"
	`include "pss_port.svh"
	`include "pss_export.svh"
endpackage

